module RISC32bitprocessor (
    input clk,
    input reset,
    input [31:0] instruction,
    output [31:0] result
);
// Your logic here
endmodule
